library verilog;
use verilog.vl_types.all;
entity booth_vlg_vec_tst is
end booth_vlg_vec_tst;
